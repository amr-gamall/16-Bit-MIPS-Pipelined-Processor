`include "aluSingleB"


module(input a, input b, output s, output c);



endmodule

